module barrelShifter16 
(
	input wire [15:0] iData,
	input wire [15:0] iRotate,
	output reg [15:0] oData
);


always @(*) begin
	case (iRotate)


	endcase
end



endmodule

